library ieee;
use ieee.std_logic_1164.all;
use work.components.all;

entity TB_MIPS is
end;

architecture impl1 of TB_MIPS is
begin
end architecture;
