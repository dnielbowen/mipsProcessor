-- Control logic
