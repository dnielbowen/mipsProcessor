library ieee;
use ieee.std_logic_1164.all;

entity MIPS_IF is
    port (
        D
    );
end;
